module subBytes128 (x, y);
input [127:0] x;
output [127:0] y;
wire [31:0] x0, x1, x2, x3;
wire [31:0] y0, y1, y2, y3;

assign x0 = x[127:96];
assign x1 = x[ 95:64];
assign x2 = x[ 63:32];
assign x3 = x[ 31: 0];

subBytes32 sub0 (x0, y0);
subBytes32 sub1 (x1, y1);
subBytes32 sub2 (x2, y2);
subBytes32 sub3 (x3, y3);

assign y = {y0, y1, y2, y3};
endmodule


module subBytes32 (x, y);
input [31:0] x;
output [31:0] y;
wire [7:0] x0, x1, x2, x3;
wire [7:0] y0, y1, y2, y3;

assign x0 = x[31:24];
assign x1 = x[23:16];
assign x2 = x[15: 8];
assign x3 = x[ 7: 0];

subBytes sub0 (x0, y0);
subBytes sub1 (x1, y1);
subBytes sub2 (x2, y2);
subBytes sub3 (x3, y3);

assign y = {y0, y1, y2, y3};
endmodule


module subBytes(x, y);
input [7:0]x;
output [7:0] y;
reg [7:0] y;

always @(x) begin
    case (x)
        /*{{{*/
        8'h00:  y <= 8'b01100011;
        8'h01:  y <= 8'b01111010;
        8'h02:  y <= 8'b01110111;
        8'h03:  y <= 8'b01111011;
        8'h04:  y <= 8'b11110010;
        8'h05:  y <= 8'b01101011;
        8'h06:  y <= 8'b01101111;
        8'h07:  y <= 8'b10110101;
        8'h08:  y <= 8'b00110000;
        8'h09:  y <= 8'b00000001;
        8'h0a:  y <= 8'b01100111;
        8'h0b:  y <= 8'b00101011;
        8'h0c:  y <= 8'b11111110;
        8'h0d:  y <= 8'b11010111;
        8'h0e:  y <= 8'b10101011;
        8'h0f:  y <= 8'b01110110;
        8'h10:  y <= 8'b11001010;
        8'h11:  y <= 8'b10000010;
        8'h12:  y <= 8'b11001001;
        8'h13:  y <= 8'b01111101;
        8'h14:  y <= 8'b11111010;
        8'h15:  y <= 8'b01011001;
        8'h16:  y <= 8'b01000111;
        8'h17:  y <= 8'b11110000;
        8'h18:  y <= 8'b10101101;
        8'h19:  y <= 8'b11010100;
        8'h1a:  y <= 8'b10100010;
        8'h1b:  y <= 8'b10101111;
        8'h1c:  y <= 8'b10011100;
        8'h1d:  y <= 8'b10100100;
        8'h1e:  y <= 8'b01110010;
        8'h1f:  y <= 8'b11000000;
        8'h20:  y <= 8'b10110111;
        8'h21:  y <= 8'b11111101;
        8'h22:  y <= 8'b10010011;
        8'h23:  y <= 8'b00100110;
        8'h24:  y <= 8'b00110110;
        8'h25:  y <= 8'b00111111;
        8'h26:  y <= 8'b11110111;
        8'h27:  y <= 8'b11001100;
        8'h28:  y <= 8'b00110100;
        8'h29:  y <= 8'b10100101;
        8'h2a:  y <= 8'b11100101;
        8'h2b:  y <= 8'b11110001;
        8'h2c:  y <= 8'b01110001;
        8'h2d:  y <= 8'b11011000;
        8'h2e:  y <= 8'b00110001;
        8'h2f:  y <= 8'b00010101;
        8'h30:  y <= 8'b00000100;
        8'h31:  y <= 8'b11000111;
        8'h32:  y <= 8'b00100011;
        8'h33:  y <= 8'b11000011;
        8'h34:  y <= 8'b00011000;
        8'h35:  y <= 8'b10010110;
        8'h36:  y <= 8'b00000101;
        8'h37:  y <= 8'b10011010;
        8'h38:  y <= 8'b00000111;
        8'h39:  y <= 8'b00010010;
        8'h3a:  y <= 8'b10000000;
        8'h3b:  y <= 8'b11100010;
        8'h3c:  y <= 8'b11101011;
        8'h3d:  y <= 8'b00100111;
        8'h3e:  y <= 8'b10110010;
        8'h3f:  y <= 8'b01110101;
        8'h40:  y <= 8'b00001001;
        8'h41:  y <= 8'b10000011;
        8'h42:  y <= 8'b00101100;
        8'h43:  y <= 8'b00011010;
        8'h44:  y <= 8'b00011011;
        8'h45:  y <= 8'b01101110;
        8'h46:  y <= 8'b01011010;
        8'h47:  y <= 8'b10100000;
        8'h48:  y <= 8'b01010010;
        8'h49:  y <= 8'b00111011;
        8'h4a:  y <= 8'b11010110;
        8'h4b:  y <= 8'b10110011;
        8'h4c:  y <= 8'b00101001;
        8'h4d:  y <= 8'b11100011;
        8'h4e:  y <= 8'b00101111;
        8'h4f:  y <= 8'b10000100;
        8'h50:  y <= 8'b01010011;
        8'h51:  y <= 8'b10110001;
        8'h52:  y <= 8'b00000000;
        8'h53:  y <= 8'b11101101;
        8'h54:  y <= 8'b00100000;
        8'h55:  y <= 8'b11111100;
        8'h56:  y <= 8'b10110001;
        8'h57:  y <= 8'b01011011;
        8'h58:  y <= 8'b01101010;
        8'h59:  y <= 8'b11001011;
        8'h5a:  y <= 8'b10111110;
        8'h5b:  y <= 8'b00111001;
        8'h5c:  y <= 8'b01001010;
        8'h5d:  y <= 8'b01001100;
        8'h5e:  y <= 8'b01011000;
        8'h5f:  y <= 8'b11001111;
        8'h60:  y <= 8'b11010000;
        8'h61:  y <= 8'b11101111;
        8'h62:  y <= 8'b10101010;
        8'h63:  y <= 8'b11111011;
        8'h64:  y <= 8'b01000011;
        8'h65:  y <= 8'b01001101;
        8'h66:  y <= 8'b00110011;
        8'h67:  y <= 8'b10000101;
        8'h68:  y <= 8'b01000101;
        8'h69:  y <= 8'b11111001;
        8'h6a:  y <= 8'b00000010;
        8'h6b:  y <= 8'b01111111;
        8'h6c:  y <= 8'b01010000;
        8'h6d:  y <= 8'b00111100;
        8'h6e:  y <= 8'b10011111;
        8'h6f:  y <= 8'b10101000;
        8'h70:  y <= 8'b01010001;
        8'h71:  y <= 8'b10100011;
        8'h72:  y <= 8'b01000000;
        8'h73:  y <= 8'b10001111;
        8'h74:  y <= 8'b10010010;
        8'h75:  y <= 8'b10011101;
        8'h76:  y <= 8'b00111000;
        8'h77:  y <= 8'b11110101;
        8'h78:  y <= 8'b10111100;
        8'h79:  y <= 8'b10110110;
        8'h7a:  y <= 8'b11011010;
        8'h7b:  y <= 8'b00100001;
        8'h7c:  y <= 8'b00010000;
        8'h7d:  y <= 8'b11111110;
        8'h7e:  y <= 8'b11110011;
        8'h7f:  y <= 8'b11010010;
        8'h80:  y <= 8'b11001101;
        8'h81:  y <= 8'b00001100;
        8'h82:  y <= 8'b00010011;
        8'h83:  y <= 8'b11101100;
        8'h84:  y <= 8'b01011111;
        8'h85:  y <= 8'b10010111;
        8'h86:  y <= 8'b01000100;
        8'h87:  y <= 8'b00010111;
        8'h88:  y <= 8'b11000100;
        8'h89:  y <= 8'b10100111;
        8'h8a:  y <= 8'b01111110;
        8'h8b:  y <= 8'b00111101;
        8'h8c:  y <= 8'b01100100;
        8'h8d:  y <= 8'b01011101;
        8'h8e:  y <= 8'b00011001;
        8'h8f:  y <= 8'b01110011;
        8'h90:  y <= 8'b01100000;
        8'h91:  y <= 8'b10000001;
        8'h92:  y <= 8'b01001111;
        8'h93:  y <= 8'b11011100;
        8'h94:  y <= 8'b00100010;
        8'h95:  y <= 8'b00101010;
        8'h96:  y <= 8'b10010000;
        8'h97:  y <= 8'b10001000;
        8'h98:  y <= 8'b01000110;
        8'h99:  y <= 8'b11101110;
        8'h9a:  y <= 8'b10111000;
        8'h9b:  y <= 8'b00010100;
        8'h9c:  y <= 8'b11011110;
        8'h9d:  y <= 8'b01011110;
        8'h9e:  y <= 8'b00001011;
        8'h9f:  y <= 8'b11011011;
        8'ha0:  y <= 8'b11100000;
        8'ha1:  y <= 8'b00110010;
        8'ha2:  y <= 8'b00111010;
        8'ha3:  y <= 8'b00001010;
        8'ha4:  y <= 8'b01001001;
        8'ha5:  y <= 8'b00000110;
        8'ha6:  y <= 8'b00100100;
        8'ha7:  y <= 8'b01011100;
        8'ha8:  y <= 8'b11000010;
        8'ha9:  y <= 8'b11010011;
        8'haa:  y <= 8'b10101100;
        8'hab:  y <= 8'b01100010;
        8'hac:  y <= 8'b10010001;
        8'had:  y <= 8'b10010101;
        8'hae:  y <= 8'b11100100;
        8'haf:  y <= 8'b01111001;
        8'hb0:  y <= 8'b11100111;
        8'hb1:  y <= 8'b11001000;
        8'hb2:  y <= 8'b00110111;
        8'hb3:  y <= 8'b01101101;
        8'hb4:  y <= 8'b10001101;
        8'hb5:  y <= 8'b11010101;
        8'hb6:  y <= 8'b01001110;
        8'hb7:  y <= 8'b10101001;
        8'hb8:  y <= 8'b01101100;
        8'hb9:  y <= 8'b01010110;
        8'hba:  y <= 8'b11110100;
        8'hbb:  y <= 8'b11101010;
        8'hbc:  y <= 8'b01100101;
        8'hbd:  y <= 8'b01111010;
        8'hbe:  y <= 8'b10101110;
        8'hbf:  y <= 8'b00001000;
        8'hc0:  y <= 8'b10111010;
        8'hc1:  y <= 8'b01111000;
        8'hc2:  y <= 8'b00100101;
        8'hc3:  y <= 8'b00101110;
        8'hc4:  y <= 8'b00011100;
        8'hc5:  y <= 8'b10100110;
        8'hc6:  y <= 8'b10110100;
        8'hc7:  y <= 8'b11000110;
        8'hc8:  y <= 8'b11101000;
        8'hc9:  y <= 8'b11011101;
        8'hca:  y <= 8'b01110100;
        8'hcb:  y <= 8'b00011111;
        8'hcc:  y <= 8'b01001011;
        8'hcd:  y <= 8'b10111101;
        8'hce:  y <= 8'b10001011;
        8'hcf:  y <= 8'b10001010;
        8'hd0:  y <= 8'b01110000;
        8'hd1:  y <= 8'b00111110;
        8'hd2:  y <= 8'b10110101;
        8'hd3:  y <= 8'b01100110;
        8'hd4:  y <= 8'b01001000;
        8'hd5:  y <= 8'b00000011;
        8'hd6:  y <= 8'b11110110;
        8'hd7:  y <= 8'b00001110;
        8'hd8:  y <= 8'b01100001;
        8'hd9:  y <= 8'b00110101;
        8'hda:  y <= 8'b01010111;
        8'hdb:  y <= 8'b10111001;
        8'hdc:  y <= 8'b10000110;
        8'hdd:  y <= 8'b11000001;
        8'hde:  y <= 8'b00011101;
        8'hdf:  y <= 8'b10011110;
        8'he0:  y <= 8'b11100001;
        8'he1:  y <= 8'b11111000;
        8'he2:  y <= 8'b10011000;
        8'he3:  y <= 8'b00010001;
        8'he4:  y <= 8'b01101001;
        8'he5:  y <= 8'b11011001;
        8'he6:  y <= 8'b10001110;
        8'he7:  y <= 8'b10010100;
        8'he8:  y <= 8'b10011011;
        8'he9:  y <= 8'b00011110;
        8'hea:  y <= 8'b10000111;
        8'heb:  y <= 8'b11101001;
        8'hec:  y <= 8'b11001110;
        8'hed:  y <= 8'b01010101;
        8'hee:  y <= 8'b00101000;
        8'hef:  y <= 8'b11011111;
        8'hf0:  y <= 8'b10001100;
        8'hf1:  y <= 8'b10100001;
        8'hf2:  y <= 8'b10001001;
        8'hf3:  y <= 8'b00001101;
        8'hf4:  y <= 8'b10111111;
        8'hf5:  y <= 8'b11100110;
        8'hf6:  y <= 8'b01000010;
        8'hf7:  y <= 8'b01101000;
        8'hf8:  y <= 8'b01000001;
        8'hf9:  y <= 8'b10011001;
        8'hfa:  y <= 8'b00101101;
        8'hfb:  y <= 8'b00001111;
        8'hfc:  y <= 8'b10110000;
        8'hfd:  y <= 8'b01010100;
        8'hfe:  y <= 8'b10111011;
        8'hff:  y <= 8'b00010110;/*}}}*/
    endcase
end
endmodule
