module expandKey_inv (in, count, out);
input [127:0] in;
input [7:0] count;
output [127:0] out;
wire [31:0] in0, in1, in2, in3;
wire [31:0] out0, out1, out2, out3;
wire [31:0] rc, rw, sw, rt;
wire [7:0]cot;
assign cot = 8'h14 - count;
assign in0 = in[127:96];
assign in1 = in[ 95:64];
assign in2 = in[ 63:32];
assign in3 = in[ 31: 0];
assign out3 = in2 ^ in3;
assign out2 = in2 ^ in1;
assign out1 = in1 ^ in0;
assign rw = (out3 & 32'hff000000) >> 24 | (out3 & 32'h00ffffff) << 8;
subBytes32 sub (rw, sw);
assign rc = (cot > 8'h08)? (32'h1b000000 << (cot - 8'h09)) : (32'h01000000 << (cot - 1));
assign rt = sw ^ rc;
assign out0 = in0 ^ rt;
assign out = {out0, out1, out2, out3};
endmodule
