module Trivium_Comp (Kin,       //IN  80bit   KEY  input
                     Din,       //IN  80bit   IV   input
                     Dout,      //OUT 512Byte Date output
                     Krdy,      //IN  1bit
                     Drdy,      //IN  1bit
                     EncDec,    //IN  1bit    1->decryption, 0->encription
                     RSTn,      //IN  1bit    reset
                     EN,        //IN  1bit    enable
                     CLK,       //IN  1bit    clk
                     BSY,       //OUT 1bit    encription or decryption time
                     Kvld,      //OUT 1bit    key generation complete
                     Dvld);     //OUT 1bit    encription or decryption complete

// input [159:0]  Kin;
// input [4095:0] Din;
input [79:0] Kin;
input [79:0] Din;
input Krey, Drdy, EncDec, RSTn, EN, CLK;
output [4095:0] Dout;
output BSY, Kvld, Dvld;

wire [15:0] fst, max;
wire [79:0] li_iv, li_key;
reg [15:0] count;
reg [287:0] SET;
reg t1, t2, t3;
reg BSYrg, Kvldrg, Dvkdrg;
reg [4095:0] z;

assign len = 4095;
assign fst = 1152;
assign max = fst + len;
assign li_key = {Kin[7:0],   Kin[15:8],  Kin[23:16],  Kin[31:24],   Kin[39:32],   Kin[47:40],   Kin[55:48],   Kin[63:56],   Kin[71:64],   Kin[79:72]};
assign li_iv  = {Din[7:0],   Din[15:8],  Din[23:16],  Din[31:24],   Din[39:32],   Din[47:40],   Din[55:48],   Din[63:56],   Din[71:64],   Din[79:72]};
// assign li_iv  = {Kin[87:80], Kin[95:88], Kin[103:96], Kin[111:104], Kin[119:112], Kin[127:120], Kin[135:128], Kin[143:136], Kin[151:144], Kin[159:152]};

always @(posedge CLK) begin
    if(RSTn == 0) begin
        SET    <= 0;
        count  <= 0;
        BSYrg  <= 0;
        Kvldrg <= 0;
        Dvldrg <= 0;
    end else if(EN == 1) begin
        if(EncDec) begin
            if(Krdy) begin
                SET   <= {3'b111, 112'b0, li_iv, 13'b0, li_key};
                count <= count + 1;
                assign Kvld = 1;
            end else begin
            end
            if(count < max) begin
                if(count == 0) begin
                end
                t1 = SET[65]  ^ SET[92];
                t2 = SET[161] ^ SET[176];
                t3 = SET[242] ^ SET[287];
                if(fst <= count) begin
                    z[len - count + fst - 1] = t1 ^ t2 ^ t3;
                end
                t1 = t1 ^ (SET[90]  & SET[91] ) ^ SET[170];
                t2 = t2 ^ (SET[174] & SET[175]) ^ SET[263];
                t3 = t3 ^ (SET[285] & SET[286]) ^ SET[68];
                SET   <= {SET[286:177], t2, SET[175:93], t1, SET[91:0], t3};
                count <= count + 1;
            end else begin
                re_OUT <= z;
            end
        end
    end
end

endmodule

