module roundFunc (word, key, count, roundWord);
    input [127:0] word;
    input [7:0] count;
    output [127:0] roundWord;
endmodule
