module test;
    
endmodule
