// and_2
module and_2 (IN1, IN2, OUT);
    input IN1, IN2;
    output OUT;
    and U1 (OUT, IN1, IN2);
endmodule
